module top_module ( input a, input b, output out );
    mod_a ins1(a,b,out);
endmodule